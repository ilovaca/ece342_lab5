module LDA_peripheral ();


endmodule
